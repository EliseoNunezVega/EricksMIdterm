`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/26/2016 07:38:27 PM
// Design Name: 
// Module Name: 1bit_alu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module 1bit_alu(
    input op1,
    input op2,
    input opsel,
    input node,
    output result,
    output c_flag,
    output z_flag,
    output o_flag,
    output s_flag
    );
endmodule
